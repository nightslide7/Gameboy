module mmio(/*AUTOARG*/);
   
endmodule
